// Demonstrate Auto-Connect features

module DffTester(input in, out);

output out;
reg out;


endmodule
