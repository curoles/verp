// // Demonstrate Auto-Connect /*features*/

/* module DffTester
 *
 */
module DffTester(input in, out);

output out;;;
reg out;

aa = bbb+cc;

endmodule
