// // Demonstrate Auto-Connect /*features*/

/* module DffTester
 *
 */
module DffTester(input in, out);

output out;;;
reg out;

aa = bbb+cc;

endmodule

  /*s o me other module*/
module 
Test2(a, output b);

endmodule
